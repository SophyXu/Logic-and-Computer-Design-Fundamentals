module shift_reg(clk, S, s_in, p_in, Q);
input wire clk, S, s_in;
input wire [15:0] p_in;
output wire [15:0] Q;
wire D[15:0];
wire nS;
FD FDQ0(.C(clk), .D(D[0]), .Q(Q[0])),
FDQ1(.C(clk), .D(D[1]), .Q(Q[1])),
FDQ2(.C(clk), .D(D[2]), .Q(Q[2])),
FDQ3(.C(clk), .D(D[3]), .Q(Q[3])),
FDQ4(.C(clk), .D(D[4]), .Q(Q[4])),
FDQ5(.C(clk), .D(D[5]), .Q(Q[5])), 
FDQ6(.C(clk), .D(D[6]), .Q(Q[6])),
FDQ7(.C(clk), .D(D[7]), .Q(Q[7])),
FDQ8(.C(clk), .D(D[8]), .Q(Q[8])),
FDQ9(.C(clk), .D(D[9]), .Q(Q[9])),
FDQ10(.C(clk), .D(D[10]), .Q(Q[10])),
FDQ11(.C(clk), .D(D[11]), .Q(Q[11])),
FDQ12(.C(clk), .D(D[12]), .Q(Q[12])),
FDQ13(.C(clk), .D(D[13]), .Q(Q[13])),
FDQ14(.C(clk), .D(D[14]), .Q(Q[14])),
FDQ15(.C(clk), .D(D[15]), .Q(Q[15]));
OR2 D0_L(.I0(L_0), .I1(R_0), .O(D[0])), 
D1_L(.I0(L_1), .I1(R_1), .O(D[1])),
D2_L(.I0(L_2), .I1(R_2), .O(D[2])),
D3_L(.I0(L_3), .I1(R_3), .O(D[3])),
D4_L(.I0(L_4), .I1(R_4), .O(D[4])),
D5_L(.I0(L_5), .I1(R_5), .O(D[5])),
D6_L(.I0(L_6), .I1(R_6), .O(D[6])),
D7_L(.I0(L_7), .I1(R_7), .O(D[7])),
D8_L(.I0(L_8), .I1(R_8), .O(D[8])),
D9_L(.I0(L_9), .I1(R_9), .O(D[9])),
D10_L(.I0(L_10), .I1(R_10), .O(D[10])),
D11_L(.I0(L_11), .I1(R_11), .O(D[11])),
D12_L(.I0(L_12), .I1(R_12), .O(D[12])),
D13_L(.I0(L_13), .I1(R_13), .O(D[13])),
D14_L(.I0(L_14), .I1(R_14), .O(D[14])),
D15_L(.I0(L_15), .I1(R_15), .O(D[15]));
AND2 L0_L(.I0(Q[1]), .I1(nS), .O(L_0)), 
L1_L(.I0(Q[2]), .I1(nS), .O(L_1)),
L2_L(.I0(Q[3]), .I1(nS), .O(L_2)),
L3_L(.I0(Q[4]), .I1(nS), .O(L_3)),
L4_L(.I0(Q[5]), .I1(nS), .O(L_4)),
L5_L(.I0(Q[6]), .I1(nS), .O(L_5)),
L6_L(.I0(Q[7]), .I1(nS), .O(L_6)),
L7_L(.I0(Q[8]), .I1(nS), .O(L_7)),
L8_L(.I0(Q[9]), .I1(nS), .O(L_8)),
L9_L(.I0(Q[10]), .I1(nS), .O(L_9)),
L10_L(.I0(Q[11]), .I1(nS), .O(L_10)),
L11_L(.I0(Q[12]), .I1(nS), .O(L_11)),
L12_L(.I0(Q[13]), .I1(nS), .O(L_12)),
L13_L(.I0(Q[14]), .I1(nS), .O(L_13)),
L14_L(.I0(Q[15]), .I1(nS), .O(L_14)),
L15_L(.I0(s_in), .I1(nS), .O(L_15));
AND2 R0_L(.I0(p_in[0]), .I1(S), .O(R_0)), 
R1_L(.I0(p_in[1]), .I1(S), .O(R_1)),
R2_L(.I0(p_in[2]), .I1(S), .O(R_2)),
R3_L(.I0(p_in[3]), .I1(S), .O(R_3)),
R4_L(.I0(p_in[4]), .I1(S), .O(R_4)),
R5_L(.I0(p_in[5]), .I1(S), .O(R_5)),
R6_L(.I0(p_in[6]), .I1(S), .O(R_6)),
R7_L(.I0(p_in[7]), .I1(S), .O(R_7)),
R8_L(.I0(p_in[8]), .I1(S), .O(R_8)),
R9_L(.I0(p_in[9]), .I1(S), .O(R_9)),
R10_L(.I0(p_in[10]), .I1(S), .O(R_10)),
R11_L(.I0(p_in[11]), .I1(S), .O(R_11)),
R12_L(.I0(p_in[12]), .I1(S), .O(R_12)),
R13_L(.I0(p_in[13]), .I1(S), .O(R_13)),
R14_L(.I0(p_in[14]), .I1(S), .O(R_14)),
R15_L(.I0(p_in[15]), .I1(S), .O(R_15));
INV nS_L(.I(S), .O(nS));
endmodule 

